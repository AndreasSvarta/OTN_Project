library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
use std.textio.all;

entity frm_scramble is
port (
	clk	: in std_logic;
	rst	: in std_logic;
	in_dat	: in std_logic_vector(255 downto 0);
	in_val	: in std_logic;
	out_val	: out std_logic;
	row	: in std_logic_vector(1 downto 0);
	column : in std_logic_vector(6 downto 0);
	out_dat	: out std_logic_vector(255 downto 0)
	);
end entity;


architecture frm_scramble_arch of frm_scramble is

signal out_dat_temp      : std_logic_vector(255 downto 0) :=(others => '0');
signal s_reg	         : std_logic_vector(15 downto 0)  :="1111111111111111";
constant s_reg_init : std_logic_vector(15 downto 0) := "1111111111111111";

begin


process (clk)
begin
if (rising_edge(clk)) then 
if (column = "0000000" and row = "00") then

out_dat_temp(255) <= in_dat(255);
out_dat_temp(254) <= in_dat(254);
out_dat_temp(253) <= in_dat(253);
out_dat_temp(252) <= in_dat(252);
out_dat_temp(251) <= in_dat(251);
out_dat_temp(250) <= in_dat(250);
out_dat_temp(249) <= in_dat(249);
out_dat_temp(248) <= in_dat(248);
out_dat_temp(247) <= in_dat(247);
out_dat_temp(246) <= in_dat(246);
out_dat_temp(245) <= in_dat(245);
out_dat_temp(244) <= in_dat(244);
out_dat_temp(243) <= in_dat(243);
out_dat_temp(242) <= in_dat(242);
out_dat_temp(241) <= in_dat(241);
out_dat_temp(240) <= in_dat(240);
out_dat_temp(239) <= in_dat(239);
out_dat_temp(238) <= in_dat(238);
out_dat_temp(237) <= in_dat(237);
out_dat_temp(236) <= in_dat(236);
out_dat_temp(235) <= in_dat(235);
out_dat_temp(234) <= in_dat(234);
out_dat_temp(233) <= in_dat(233);
out_dat_temp(232) <= in_dat(232);
out_dat_temp(231) <= in_dat(231);
out_dat_temp(230) <= in_dat(230);
out_dat_temp(229) <= in_dat(229);
out_dat_temp(228) <= in_dat(228);
out_dat_temp(227) <= in_dat(227);
out_dat_temp(226) <= in_dat(226);
out_dat_temp(225) <= in_dat(225);
out_dat_temp(224) <= in_dat(224);
out_dat_temp(223) <= in_dat(223);
out_dat_temp(222) <= in_dat(222);
out_dat_temp(221) <= in_dat(221);
out_dat_temp(220) <= in_dat(220);
out_dat_temp(219) <= in_dat(219);
out_dat_temp(218) <= in_dat(218);
out_dat_temp(217) <= in_dat(217);
out_dat_temp(216) <= in_dat(216);
out_dat_temp(215) <= in_dat(215);
out_dat_temp(214) <= in_dat(214);
out_dat_temp(213) <= in_dat(213);
out_dat_temp(212) <= in_dat(212);
out_dat_temp(211) <= in_dat(211);
out_dat_temp(210) <= in_dat(210);
out_dat_temp(209) <= in_dat(209);
out_dat_temp(208) <= in_dat(208);
out_dat_temp(207)  <= in_dat(207) xor s_reg_init(15);
out_dat_temp(206)  <= in_dat(206) xor s_reg_init(14);
out_dat_temp(205)  <= in_dat(205) xor s_reg_init(13);
out_dat_temp(204)  <= in_dat(204) xor s_reg_init(12);
out_dat_temp(203)  <= in_dat(203) xor s_reg_init(11);
out_dat_temp(202)  <= in_dat(202) xor s_reg_init(10);
out_dat_temp(201)  <= in_dat(201) xor s_reg_init(9);
out_dat_temp(200)  <= in_dat(200) xor s_reg_init(8);
out_dat_temp(199)  <= in_dat(199) xor s_reg_init(7);
out_dat_temp(198)  <= in_dat(198) xor s_reg_init(6);
out_dat_temp(197)  <= in_dat(197) xor s_reg_init(5);
out_dat_temp(196)  <= in_dat(196) xor s_reg_init(4);
out_dat_temp(195)  <= in_dat(195) xor s_reg_init(3);
out_dat_temp(194)  <= in_dat(194) xor s_reg_init(2);
out_dat_temp(193)  <= in_dat(193) xor s_reg_init(1);
out_dat_temp(192)  <= in_dat(192) xor s_reg_init(0);
out_dat_temp(191)  <= in_dat(191) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(190)  <= in_dat(190) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(189)  <= in_dat(189) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(188)  <= in_dat(188) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(187)  <= in_dat(187) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(2);
out_dat_temp(186)  <= in_dat(186) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(1);
out_dat_temp(185)  <= in_dat(185) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(0);
out_dat_temp(184)  <= in_dat(184) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(183)  <= in_dat(183) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(182)  <= in_dat(182) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(181)  <= in_dat(181) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(180)  <= in_dat(180) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(179)  <= in_dat(179) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(178)  <= in_dat(178) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(177)  <= in_dat(177) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(176)  <= in_dat(176) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(175)  <= in_dat(175) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(8) xor s_reg_init(4);
out_dat_temp(174)  <= in_dat(174) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(7) xor s_reg_init(3);
out_dat_temp(173)  <= in_dat(173) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(6) xor s_reg_init(2);
out_dat_temp(172)  <= in_dat(172) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(5) xor s_reg_init(1);
out_dat_temp(171)  <= in_dat(171) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(4) xor s_reg_init(0);
out_dat_temp(170)  <= in_dat(170) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(169)  <= in_dat(169) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(168)  <= in_dat(168) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(2);
out_dat_temp(167)  <= in_dat(167) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(1);
out_dat_temp(166)  <= in_dat(166) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(0);
out_dat_temp(165)  <= in_dat(165) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(164)  <= in_dat(164) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(163)  <= in_dat(163) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(162)  <= in_dat(162) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(161)  <= in_dat(161) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(160)  <= in_dat(160) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(3);
out_dat_temp(159)  <= in_dat(159) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(158)  <= in_dat(158) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(157)  <= in_dat(157) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(156)  <= in_dat(156)xor s_reg_init(15) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(155)  <= in_dat(155) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(154)  <= in_dat(154) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(153)  <= in_dat(153) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(152)  <= in_dat(152) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(151)  <= in_dat(151) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(150)  <= in_dat(150) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(149)  <= in_dat(149) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(148)  <= in_dat(148) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4);
out_dat_temp(147)  <= in_dat(147) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3);
out_dat_temp(146)  <= in_dat(146) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(145)  <= in_dat(145) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(144)  <= in_dat(144) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(143)  <= in_dat(143) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(142)  <= in_dat(142) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(141)  <= in_dat(141) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(140)  <= in_dat(140) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(139)  <= in_dat(139) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(138)  <= in_dat(138) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5);
out_dat_temp(137)  <= in_dat(137) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4);
out_dat_temp(136)  <= in_dat(136) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3);
out_dat_temp(135)  <= in_dat(135) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(134)  <= in_dat(134) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(133)  <= in_dat(133) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(132)  <= in_dat(132) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(131)  <= in_dat(131) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(130)  <= in_dat(130) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(2);
out_dat_temp(129)  <= in_dat(129) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(1);
out_dat_temp(128)  <= in_dat(128) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(0);
out_dat_temp(127)  <= in_dat(127) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(126)  <= in_dat(126) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(125)  <= in_dat(125) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4);
out_dat_temp(124)  <= in_dat(124) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3);
out_dat_temp(123)  <= in_dat(123) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(122)  <= in_dat(122) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(121)  <= in_dat(121) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(120)  <= in_dat(120) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(119)  <= in_dat(119) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(118)  <= in_dat(118) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(117)  <= in_dat(117) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(116)  <= in_dat(116) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(1);
out_dat_temp(115)  <= in_dat(115) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(0);
out_dat_temp(114)  <= in_dat(114) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(0);
out_dat_temp(113)  <= in_dat(113) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(0);
out_dat_temp(112)  <= in_dat(112) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(0);
out_dat_temp(111)  <= in_dat(111) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(0);
out_dat_temp(110)  <= in_dat(110) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(0);
out_dat_temp(109)  <= in_dat(109) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(108)  <= in_dat(108) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(107)  <= in_dat(107) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(106)  <= in_dat(106) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(105)  <= in_dat(105) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(104)  <= in_dat(104) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(103)  <= in_dat(103) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(102)  <= in_dat(102) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7);
out_dat_temp(101)  <= in_dat(101) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6);
out_dat_temp(100)  <= in_dat(100) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5);
out_dat_temp(99)  <= in_dat(99) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4);
out_dat_temp(98)  <= in_dat(98) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3);
out_dat_temp(97)  <= in_dat(97) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(96)  <= in_dat(96) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(95)  <= in_dat(95) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(94)  <= in_dat(94) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3);
out_dat_temp(93)  <= in_dat(93) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(92)  <= in_dat(92) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(91)  <= in_dat(91) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(90)  <= in_dat(90) xor s_reg_init(15) xor s_reg_init(7) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(89)  <= in_dat(89) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(6) xor s_reg_init(1);
out_dat_temp(88)  <= in_dat(88) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(5) xor s_reg_init(0);
out_dat_temp(87)  <= in_dat(87) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(86)  <= in_dat(86) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(85)  <= in_dat(85) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(1);
out_dat_temp(84)  <= in_dat(84) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(0);
out_dat_temp(83)  <= in_dat(83) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(82)  <= in_dat(82) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(81)  <= in_dat(81) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(80)  <= in_dat(80) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(79)  <= in_dat(79) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(78)  <= in_dat(78) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(77)  <= in_dat(77) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(76)  <= in_dat(76) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(75)  <= in_dat(75) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(8) xor s_reg_init(2);
out_dat_temp(74)  <= in_dat(74) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(7) xor s_reg_init(1);
out_dat_temp(73)  <= in_dat(73) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(6) xor s_reg_init(0);
out_dat_temp(72)  <= in_dat(72) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(71)  <= in_dat(71) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(70)  <= in_dat(70) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(69)  <= in_dat(69) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(68)  <= in_dat(68) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(67)  <= in_dat(67) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(66)  <= in_dat(66) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(65)  <= in_dat(65) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(64)  <= in_dat(64) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(63)  <= in_dat(63) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(62)  <= in_dat(62) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(61)  <= in_dat(61) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(60)  <= in_dat(60) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(59)  <= in_dat(59) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(58)  <= in_dat(58) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(57)  <= in_dat(57) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(56)  <= in_dat(56) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(55)  <= in_dat(55) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(54)  <= in_dat(54) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(53)  <= in_dat(53) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(52)  <= in_dat(52) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(51)  <= in_dat(51) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(50)  <= in_dat(50) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(49)  <= in_dat(49) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(48)  <= in_dat(48) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(47)  <= in_dat(47) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(46)  <= in_dat(46) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(45)  <= in_dat(45) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(44)  <= in_dat(44) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(43)  <= in_dat(43) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(42)  <= in_dat(42) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(41)  <= in_dat(41) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(40)  <= in_dat(40) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(39)  <= in_dat(39) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(38)  <= in_dat(38) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(37)  <= in_dat(37) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(36)  <= in_dat(36) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4);
out_dat_temp(35)  <= in_dat(35) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3);
out_dat_temp(34)  <= in_dat(34) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(33)  <= in_dat(33) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(32)  <= in_dat(32) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(31)  <= in_dat(31) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(5);
out_dat_temp(30)  <= in_dat(30) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(4);
out_dat_temp(29)  <= in_dat(29) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(3);
out_dat_temp(28)  <= in_dat(28) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(27)  <= in_dat(27) xor s_reg_init(11) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(26)  <= in_dat(26) xor s_reg_init(10) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(25)  <= in_dat(25) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(5) xor s_reg_init(4);
out_dat_temp(24)  <= in_dat(24) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(4) xor s_reg_init(3);
out_dat_temp(23)  <= in_dat(23) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(3) xor s_reg_init(2);
out_dat_temp(22)  <= in_dat(22) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(21)  <= in_dat(21) xor s_reg_init(11) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(20)  <= in_dat(20) xor s_reg_init(15) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2);
out_dat_temp(19)  <= in_dat(19) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(18)  <= in_dat(18) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(17)  <= in_dat(17) xor s_reg_init(15) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(16)  <= in_dat(16) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(1);
out_dat_temp(15)  <= in_dat(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(0);
out_dat_temp(14)  <= in_dat(14) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(13)  <= in_dat(13) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(12)  <= in_dat(12) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(1);
out_dat_temp(11)  <= in_dat(11) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(0);
out_dat_temp(10)  <= in_dat(10) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(9)  <= in_dat(9) xor s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(8)  <= in_dat(8) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(7)  <= in_dat(7) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
out_dat_temp(6)  <= in_dat(6) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
out_dat_temp(5)  <= in_dat(5) xor s_reg_init(15) xor s_reg_init(13) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8);
out_dat_temp(4)  <= in_dat(4) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7);
out_dat_temp(3)  <= in_dat(3) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6);
out_dat_temp(2)  <= in_dat(2) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5);
out_dat_temp(1)  <= in_dat(1) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(4);
out_dat_temp(0)  <= in_dat(0) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(5) xor s_reg_init(4) xor s_reg_init(3);


s_reg(15) <= s_reg_init(9) xor s_reg_init(7) xor s_reg_init(4) xor s_reg_init(3) xor s_reg_init(2);
s_reg(14) <= s_reg_init(8) xor s_reg_init(6) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1);
s_reg(13) <= s_reg_init(7) xor s_reg_init(5) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
s_reg(12) <= s_reg_init(15) xor s_reg_init(11) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(1);
s_reg(11) <= s_reg_init(14) xor s_reg_init(10) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(1) xor s_reg_init(0);
s_reg(10) <= s_reg_init(15) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(4);
s_reg(9) <= s_reg_init(14) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(3);
s_reg(8) <= s_reg_init(13) xor s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(2);
s_reg(7) <= s_reg_init(12) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(1);
s_reg(6) <= s_reg_init(11) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(0);
s_reg(5) <= s_reg_init(15) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(2) xor s_reg_init(0);
s_reg(4) <= s_reg_init(15) xor s_reg_init(14) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(1) xor s_reg_init(0);
s_reg(3) <= s_reg_init(15) xor s_reg_init(14) xor s_reg_init(13) xor s_reg_init(11) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(1);
s_reg(2) <= s_reg_init(14) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(10) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(0);
s_reg(1) <= s_reg_init(15) xor s_reg_init(13) xor s_reg_init(12) xor s_reg_init(9) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(4) xor s_reg_init(0);
s_reg(0) <= s_reg_init(15) xor s_reg_init(14) xor s_reg_init(12) xor s_reg_init(8) xor s_reg_init(7) xor s_reg_init(6) xor s_reg_init(5) xor s_reg_init(3) xor s_reg_init(2) xor s_reg_init(0);


else

out_dat_temp(255)<=in_dat(255) xor s_reg(15) ;
out_dat_temp(254)<=in_dat(254) xor s_reg(14) ;
out_dat_temp(253)<=in_dat(253) xor s_reg(13) ;
out_dat_temp(252)<=in_dat(252) xor s_reg(12) ;
out_dat_temp(251)<=in_dat(251) xor s_reg(11) ;
out_dat_temp(250)<=in_dat(250) xor s_reg(10) ;
out_dat_temp(249)<=in_dat(249) xor s_reg(9) ;
out_dat_temp(248)<=in_dat(248) xor s_reg(8) ;
out_dat_temp(247)<=in_dat(247) xor s_reg(7) ;
out_dat_temp(246)<=in_dat(246) xor s_reg(6) ;
out_dat_temp(245)<=in_dat(245) xor s_reg(5) ;
out_dat_temp(244)<=in_dat(244) xor s_reg(4) ;
out_dat_temp(243)<=in_dat(243) xor s_reg(3) ;
out_dat_temp(242)<=in_dat(242) xor s_reg(2) ;
out_dat_temp(241)<=in_dat(241) xor s_reg(1) ;
out_dat_temp(240)<=in_dat(240) xor s_reg(0) ;
out_dat_temp(239)<=in_dat(239) xor s_reg(15) xor s_reg(11) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(238)<=in_dat(238) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(237)<=in_dat(237) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(236)<=in_dat(236) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(235)<=in_dat(235) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(2) ;
out_dat_temp(234)<=in_dat(234) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(1) ;
out_dat_temp(233)<=in_dat(233) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(0) ;
out_dat_temp(232)<=in_dat(232) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(231)<=in_dat(231) xor s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(230)<=in_dat(230) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(229)<=in_dat(229) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(228)<=in_dat(228) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(227)<=in_dat(227) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(226)<=in_dat(226) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(225)<=in_dat(225) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(224)<=in_dat(224) xor s_reg(15) xor s_reg(12) xor s_reg(9) xor s_reg(5) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(223)<=in_dat(223) xor s_reg(15) xor s_reg(14) xor s_reg(8) xor s_reg(4) ;
out_dat_temp(222)<=in_dat(222) xor s_reg(14) xor s_reg(13) xor s_reg(7) xor s_reg(3) ;
out_dat_temp(221)<=in_dat(221) xor s_reg(13) xor s_reg(12) xor s_reg(6) xor s_reg(2) ;
out_dat_temp(220)<=in_dat(220) xor s_reg(12) xor s_reg(11) xor s_reg(5) xor s_reg(1) ;
out_dat_temp(219)<=in_dat(219) xor s_reg(11) xor s_reg(10) xor s_reg(4) xor s_reg(0) ;
out_dat_temp(218)<=in_dat(218) xor s_reg(15) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(217)<=in_dat(217) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(216)<=in_dat(216) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(2) ;
out_dat_temp(215)<=in_dat(215) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(1) ;
out_dat_temp(214)<=in_dat(214) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(0) ;
out_dat_temp(213)<=in_dat(213) xor s_reg(15) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(212)<=in_dat(212) xor s_reg(15) xor s_reg(14) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(211)<=in_dat(211) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(210)<=in_dat(210) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(209)<=in_dat(209) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(208)<=in_dat(208) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(8) xor s_reg(5) xor s_reg(3) ;
out_dat_temp(207)<=in_dat(207) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(7) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(206)<=in_dat(206) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(6) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(205)<=in_dat(205) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(5) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(204)<=in_dat(204) xor s_reg(15) xor s_reg(10) xor s_reg(8) xor s_reg(4) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(203)<=in_dat(203) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(202)<=in_dat(202) xor s_reg(14) xor s_reg(13) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(201)<=in_dat(201) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(200)<=in_dat(200) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(199)<=in_dat(199) xor s_reg(15) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(198)<=in_dat(198) xor s_reg(14) xor s_reg(12) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(197)<=in_dat(197) xor s_reg(13) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(196)<=in_dat(196) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(4) ;
out_dat_temp(195)<=in_dat(195) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(3) ;
out_dat_temp(194)<=in_dat(194) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(193)<=in_dat(193) xor s_reg(12) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(192)<=in_dat(192) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(191)<=in_dat(191) xor s_reg(15) xor s_reg(11) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(190)<=in_dat(190) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(189)<=in_dat(189) xor s_reg(14) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(188)<=in_dat(188) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(187)<=in_dat(187) xor s_reg(15) xor s_reg(12) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(186)<=in_dat(186) xor s_reg(15) xor s_reg(14) xor s_reg(7) xor s_reg(6) xor s_reg(5) ;
out_dat_temp(185)<=in_dat(185) xor s_reg(14) xor s_reg(13) xor s_reg(6) xor s_reg(5) xor s_reg(4) ;
out_dat_temp(184)<=in_dat(184) xor s_reg(13) xor s_reg(12) xor s_reg(5) xor s_reg(4) xor s_reg(3) ;
out_dat_temp(183)<=in_dat(183) xor s_reg(12) xor s_reg(11) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(182)<=in_dat(182) xor s_reg(11) xor s_reg(10) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(181)<=in_dat(181) xor s_reg(10) xor s_reg(9) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(180)<=in_dat(180) xor s_reg(15) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(179)<=in_dat(179) xor s_reg(14) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(178)<=in_dat(178) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(2) ;
out_dat_temp(177)<=in_dat(177) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(1) ;
out_dat_temp(176)<=in_dat(176) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(0) ;
out_dat_temp(175)<=in_dat(175) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(174)<=in_dat(174) xor s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(173)<=in_dat(173) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(4) ;
out_dat_temp(172)<=in_dat(172) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(3) ;
out_dat_temp(171)<=in_dat(171) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(170)<=in_dat(170) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(169)<=in_dat(169) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(168)<=in_dat(168) xor s_reg(15) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(167)<=in_dat(167) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(166)<=in_dat(166) xor s_reg(14) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(165)<=in_dat(165) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(164)<=in_dat(164) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(1) ;
out_dat_temp(163)<=in_dat(163) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(162)<=in_dat(162) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(161)<=in_dat(161) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(160)<=in_dat(160) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(159)<=in_dat(159) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(158)<=in_dat(158) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(0) ;
out_dat_temp(157)<=in_dat(157) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(156)<=in_dat(156) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(155)<=in_dat(155) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(154)<=in_dat(154) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(153)<=in_dat(153) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(5) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(152)<=in_dat(152) xor s_reg(15) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(151)<=in_dat(151) xor s_reg(14) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(150)<=in_dat(150) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(7) ;
out_dat_temp(149)<=in_dat(149) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(6) ;
out_dat_temp(148)<=in_dat(148) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(5) ;
out_dat_temp(147)<=in_dat(147) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(4) ;
out_dat_temp(146)<=in_dat(146) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(3) ;
out_dat_temp(145)<=in_dat(145) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(144)<=in_dat(144) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(143)<=in_dat(143) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(142)<=in_dat(142) xor s_reg(15) xor s_reg(11) xor s_reg(7) xor s_reg(5) xor s_reg(3) ;
out_dat_temp(141)<=in_dat(141) xor s_reg(14) xor s_reg(10) xor s_reg(6) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(140)<=in_dat(140) xor s_reg(13) xor s_reg(9) xor s_reg(5) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(139)<=in_dat(139) xor s_reg(12) xor s_reg(8) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(138)<=in_dat(138) xor s_reg(15) xor s_reg(7) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(137)<=in_dat(137) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(6) xor s_reg(1) ;
out_dat_temp(136)<=in_dat(136) xor s_reg(14) xor s_reg(13) xor s_reg(10) xor s_reg(5) xor s_reg(0) ;
out_dat_temp(135)<=in_dat(135) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(134)<=in_dat(134) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(133)<=in_dat(133) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(9) xor s_reg(7) xor s_reg(1) ;
out_dat_temp(132)<=in_dat(132) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(8) xor s_reg(6) xor s_reg(0) ;
out_dat_temp(131)<=in_dat(131) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(7) xor s_reg(5) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(130)<=in_dat(130) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(129)<=in_dat(129) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(128)<=in_dat(128) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(4) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(127)<=in_dat(127) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(126)<=in_dat(126) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(125)<=in_dat(125) xor s_reg(15) xor s_reg(13) xor s_reg(10) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(124)<=in_dat(124) xor s_reg(14) xor s_reg(12) xor s_reg(9) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(123)<=in_dat(123) xor s_reg(15) xor s_reg(13) xor s_reg(8) xor s_reg(2) ;
out_dat_temp(122)<=in_dat(122) xor s_reg(14) xor s_reg(12) xor s_reg(7) xor s_reg(1) ;
out_dat_temp(121)<=in_dat(121) xor s_reg(13) xor s_reg(11) xor s_reg(6) xor s_reg(0) ;
out_dat_temp(120)<=in_dat(120) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(5) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(119)<=in_dat(119) xor s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(4) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(118)<=in_dat(118) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(117)<=in_dat(117) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(116)<=in_dat(116) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(115)<=in_dat(115) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(114)<=in_dat(114) xor s_reg(15) xor s_reg(13) xor s_reg(10) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(113)<=in_dat(113) xor s_reg(14) xor s_reg(12) xor s_reg(9) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(112)<=in_dat(112) xor s_reg(13) xor s_reg(11) xor s_reg(8) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(111)<=in_dat(111) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(7) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(110)<=in_dat(110) xor s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(6) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(109)<=in_dat(109) xor s_reg(14) xor s_reg(13) xor s_reg(9) xor s_reg(8) xor s_reg(5) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(108)<=in_dat(108) xor s_reg(13) xor s_reg(12) xor s_reg(8) xor s_reg(7) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(107)<=in_dat(107) xor s_reg(15) xor s_reg(12) xor s_reg(7) xor s_reg(6) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(106)<=in_dat(106) xor s_reg(14) xor s_reg(11) xor s_reg(6) xor s_reg(5) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(105)<=in_dat(105) xor s_reg(13) xor s_reg(10) xor s_reg(5) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(104)<=in_dat(104) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(103)<=in_dat(103) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(102)<=in_dat(102) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(101)<=in_dat(101) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(100)<=in_dat(100) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(99)<=in_dat(99) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(98)<=in_dat(98) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(97)<=in_dat(97) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(96)<=in_dat(96) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(95)<=in_dat(95) xor s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(94)<=in_dat(94) xor s_reg(14) xor s_reg(13) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(93)<=in_dat(93) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(92)<=in_dat(92) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(91)<=in_dat(91) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(90)<=in_dat(90) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(89)<=in_dat(89) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(88)<=in_dat(88) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(87)<=in_dat(87) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(86)<=in_dat(86) xor s_reg(15) xor s_reg(12) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(85)<=in_dat(85) xor s_reg(14) xor s_reg(11) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(84)<=in_dat(84) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(7) xor s_reg(5) xor s_reg(4) ;
out_dat_temp(83)<=in_dat(83) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(6) xor s_reg(4) xor s_reg(3) ;
out_dat_temp(82)<=in_dat(82) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(5) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(81)<=in_dat(81) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(80)<=in_dat(80) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(79)<=in_dat(79) xor s_reg(15) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(5) ;
out_dat_temp(78)<=in_dat(78) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(4) ;
out_dat_temp(77)<=in_dat(77) xor s_reg(13) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(3) ;
out_dat_temp(76)<=in_dat(76) xor s_reg(12) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(75)<=in_dat(75) xor s_reg(11) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(74)<=in_dat(74) xor s_reg(10) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(73)<=in_dat(73) xor s_reg(15) xor s_reg(11) xor s_reg(9) xor s_reg(5) xor s_reg(4) ;
out_dat_temp(72)<=in_dat(72) xor s_reg(14) xor s_reg(10) xor s_reg(8) xor s_reg(4) xor s_reg(3) ;
out_dat_temp(71)<=in_dat(71) xor s_reg(13) xor s_reg(9) xor s_reg(7) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(70)<=in_dat(70) xor s_reg(12) xor s_reg(8) xor s_reg(6) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(69)<=in_dat(69) xor s_reg(11) xor s_reg(7) xor s_reg(5) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(68)<=in_dat(68) xor s_reg(15) xor s_reg(11) xor s_reg(10) xor s_reg(6) xor s_reg(4) xor s_reg(2) ;
out_dat_temp(67)<=in_dat(67) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(5) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(66)<=in_dat(66) xor s_reg(13) xor s_reg(9) xor s_reg(8) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(65)<=in_dat(65) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(64)<=in_dat(64) xor s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(1) ;
out_dat_temp(63)<=in_dat(63) xor s_reg(14) xor s_reg(13) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(0) ;
out_dat_temp(62)<=in_dat(62) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(61)<=in_dat(61) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(60)<=in_dat(60) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(9) xor s_reg(6) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(59)<=in_dat(59) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(8) xor s_reg(5) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(58)<=in_dat(58) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(7) xor s_reg(4) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(57)<=in_dat(57) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(56)<=in_dat(56) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(5) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(55)<=in_dat(55) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(54)<=in_dat(54) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(53)<=in_dat(53) xor s_reg(15) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(8) ;
out_dat_temp(52)<=in_dat(52) xor s_reg(14) xor s_reg(12) xor s_reg(9) xor s_reg(8) xor s_reg(7) ;
out_dat_temp(51)<=in_dat(51) xor s_reg(13) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(6) ;
out_dat_temp(50)<=in_dat(50) xor s_reg(12) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(5) ;
out_dat_temp(49)<=in_dat(49) xor s_reg(11) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(4) ;
out_dat_temp(48)<=in_dat(48) xor s_reg(10) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(3) ;
out_dat_temp(47)<=in_dat(47) xor s_reg(9) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(46)<=in_dat(46) xor s_reg(8) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(45)<=in_dat(45) xor s_reg(7) xor s_reg(5) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(44)<=in_dat(44) xor s_reg(15) xor s_reg(11) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(43)<=in_dat(43) xor s_reg(14) xor s_reg(10) xor s_reg(5) xor s_reg(3) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(42)<=in_dat(42) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(4) ;
out_dat_temp(41)<=in_dat(41) xor s_reg(14) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(3) ;
out_dat_temp(40)<=in_dat(40) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(2) ;
out_dat_temp(39)<=in_dat(39) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(1) ;
out_dat_temp(38)<=in_dat(38) xor s_reg(11) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(0) ;
out_dat_temp(37)<=in_dat(37) xor s_reg(15) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(36)<=in_dat(36) xor s_reg(15) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(35)<=in_dat(35) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(4) xor s_reg(1) ;
out_dat_temp(34)<=in_dat(34) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(33)<=in_dat(33) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(0) ;
out_dat_temp(32)<=in_dat(32) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(31)<=in_dat(31) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(30)<=in_dat(30) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(29)<=in_dat(29) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(28)<=in_dat(28) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(27)<=in_dat(27) xor s_reg(15) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(3) xor s_reg(1) ;
out_dat_temp(26)<=in_dat(26) xor s_reg(14) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(25)<=in_dat(25) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(24)<=in_dat(24) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(23)<=in_dat(23) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(22)<=in_dat(22) xor s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) ;
out_dat_temp(21)<=in_dat(21) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(1) ;
out_dat_temp(20)<=in_dat(20) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(19)<=in_dat(19) xor s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(1) ;
out_dat_temp(18)<=in_dat(18) xor s_reg(14) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(17)<=in_dat(17) xor s_reg(15) xor s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(16)<=in_dat(16) xor s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(15)<=in_dat(15) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(14)<=in_dat(14) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(13)<=in_dat(13) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(12)<=in_dat(12) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(11)<=in_dat(11) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(10)<=in_dat(10) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(9)<=in_dat(9) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(8)<=in_dat(8) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(5) xor s_reg(3) xor s_reg(0) ;
out_dat_temp(7)<=in_dat(7) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(4) xor s_reg(0) ;
out_dat_temp(6)<=in_dat(6) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(3) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(5)<=in_dat(5) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(1) xor s_reg(0) ;
out_dat_temp(4)<=in_dat(4) xor s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(2) ;
out_dat_temp(3)<=in_dat(3) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(1) ;
out_dat_temp(2)<=in_dat(2) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(0) ;
out_dat_temp(1)<=in_dat(1) xor s_reg(15) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(2) xor s_reg(0) ;
out_dat_temp(0)<=in_dat(0) xor s_reg(15) xor s_reg(14) xor s_reg(9) xor s_reg(8) xor s_reg(2) xor s_reg(1) xor s_reg(0) ;



s_reg(15) <= s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(8) xor s_reg(7) xor s_reg(2) xor s_reg(1);
s_reg(14) <= s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(7) xor s_reg(6) xor s_reg(1) xor s_reg(0);
s_reg(13) <= s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(9) xor s_reg(6) xor s_reg(5) xor s_reg(2);
s_reg(12) <= s_reg(14) xor s_reg(12) xor s_reg(11) xor s_reg(8) xor s_reg(5) xor s_reg(4) xor s_reg(1);
s_reg(11) <= s_reg(13) xor s_reg(11) xor s_reg(10) xor s_reg(7) xor s_reg(4) xor s_reg(3) xor s_reg(0);
s_reg(10) <= s_reg(15) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(9) xor s_reg(6) xor s_reg(3) xor s_reg(0);
s_reg(9) <= s_reg(15) xor s_reg(14) xor s_reg(10) xor s_reg(9) xor s_reg(8) xor s_reg(5) xor s_reg(0);
s_reg(8) <= s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(7) xor s_reg(4) xor s_reg(2) xor s_reg(0);
s_reg(7) <= s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(6) xor s_reg(3) xor s_reg(2) xor s_reg(1) xor s_reg(0);
s_reg(6) <= s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(5) xor s_reg(1);
s_reg(5) <= s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(9) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(4) xor s_reg(0);
s_reg(4) <= s_reg(15) xor s_reg(13) xor s_reg(12) xor s_reg(10) xor s_reg(8) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(3) xor s_reg(2) xor s_reg(0);
s_reg(3) <= s_reg(15) xor s_reg(14) xor s_reg(12) xor s_reg(9) xor s_reg(7) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(1) xor s_reg(0);
s_reg(2) <= s_reg(15) xor s_reg(14) xor s_reg(13) xor s_reg(8) xor s_reg(6) xor s_reg(5) xor s_reg(3);
s_reg(1) <= s_reg(14) xor s_reg(13) xor s_reg(12) xor s_reg(7) xor s_reg(5) xor s_reg(4) xor s_reg(2);
s_reg(0) <= s_reg(13) xor s_reg(12) xor s_reg(11) xor s_reg(6) xor s_reg(4) xor s_reg(3) xor s_reg(1);




end if;
end if;

end process;


out_dat <= out_dat_temp;


end architecture;